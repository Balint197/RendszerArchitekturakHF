`timescale 1ns / 1ps
`default_nettype none

module spi_top(
    );


endmodule

`default_nettype wire