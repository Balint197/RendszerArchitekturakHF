`timescale 1ns / 1ps
`default_nettype none

module spi(
    );


endmodule

`default_nettype wire